module teste ();

endmodule 